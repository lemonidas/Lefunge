>025*"!dlrow ,olleH":v
                  v:,_@
                  >  ^

>&>~:"="-#v_$.55+,@
  ^  p41\&<      

v                               >15gv        >13gv
v           >~$&:14p13g+:15p14g`|   >:13p12g`|   >12pv
v                               >14g^        >12g^
>& 012p013p:|:                                     -1<
            >12g.25*,@

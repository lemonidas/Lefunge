055+"!dlrow ,olleH">:#,_@

v
v
v
v                 >11gv
>&~$11p&22p11g22g`|   >.25*,@
                  >22g^

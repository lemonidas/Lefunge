>&~$&+.25*,@

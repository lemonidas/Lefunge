>0&~$:#v_$.25*,@
v      <^ < 
>1-\&~$+\:^

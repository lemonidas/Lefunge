0&>:1-:v v *_$.55+,@
  ^    _$>\:^
